8 9
0 0 0
0 1 2
0 2 12
0 3 1
0 4 4
0 5 7
0 6 10
0 7 13
1 0 0
1 1 8
1 2 13
1 3 3
1 4 5
1 5 6
1 6 4
1 7 9
1 8 11
